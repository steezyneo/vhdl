module mux8to1_tb(    );

reg [7:0]I;
reg [2:0] S;
wire Y;
mux8to1 uut(I,S,Y);
initial begin
#100 I[7:0]=8'b00101101; S[2:0]=3'b000;
#100 I[7:0]=8'b00101101; S[2:0]=3'b001;
#100 I[7:0]=8'b00101101; S[2:0]=3'b010;
#100 I[7:0]=8'b00101101; S[2:0]=3'b011;
#100 I[7:0]=8'b00101101; S[2:0]=3'b100;
#100 I[7:0]=8'b00101101; S[2:0]=3'b101;
#100 I[7:0]=8'b00101101; S[2:0]=3'b110;
#100 I[7:0]=8'b00101101; S[2:0]=3'b111;
end
endmodule
